
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'hcbdc300d;
    ram_cell[       1] = 32'h0;  // 32'h7d93b8f1;
    ram_cell[       2] = 32'h0;  // 32'h3c17e6f1;
    ram_cell[       3] = 32'h0;  // 32'hfca192b0;
    ram_cell[       4] = 32'h0;  // 32'hd68fd792;
    ram_cell[       5] = 32'h0;  // 32'h255a4042;
    ram_cell[       6] = 32'h0;  // 32'h99dd4d01;
    ram_cell[       7] = 32'h0;  // 32'h41ec58d6;
    ram_cell[       8] = 32'h0;  // 32'h49df0ba5;
    ram_cell[       9] = 32'h0;  // 32'h0d9e7392;
    ram_cell[      10] = 32'h0;  // 32'h86652738;
    ram_cell[      11] = 32'h0;  // 32'h71598504;
    ram_cell[      12] = 32'h0;  // 32'h4b9ee300;
    ram_cell[      13] = 32'h0;  // 32'h5710ca28;
    ram_cell[      14] = 32'h0;  // 32'h43fe77ad;
    ram_cell[      15] = 32'h0;  // 32'hfd02622d;
    ram_cell[      16] = 32'h0;  // 32'h6cd03775;
    ram_cell[      17] = 32'h0;  // 32'hb98843cf;
    ram_cell[      18] = 32'h0;  // 32'h0a943465;
    ram_cell[      19] = 32'h0;  // 32'hd812b80b;
    ram_cell[      20] = 32'h0;  // 32'h4f40f0d0;
    ram_cell[      21] = 32'h0;  // 32'hae45842e;
    ram_cell[      22] = 32'h0;  // 32'hf72481a7;
    ram_cell[      23] = 32'h0;  // 32'h41c8071b;
    ram_cell[      24] = 32'h0;  // 32'h44f18b72;
    ram_cell[      25] = 32'h0;  // 32'hed4b7199;
    ram_cell[      26] = 32'h0;  // 32'hfb5f2d55;
    ram_cell[      27] = 32'h0;  // 32'h3fbc12ac;
    ram_cell[      28] = 32'h0;  // 32'hb7d87a6f;
    ram_cell[      29] = 32'h0;  // 32'hb7c28cd8;
    ram_cell[      30] = 32'h0;  // 32'h9b4eb8d9;
    ram_cell[      31] = 32'h0;  // 32'hb3e88420;
    ram_cell[      32] = 32'h0;  // 32'h8d37e3fb;
    ram_cell[      33] = 32'h0;  // 32'hc840b93b;
    ram_cell[      34] = 32'h0;  // 32'h084129a4;
    ram_cell[      35] = 32'h0;  // 32'h7ddbd766;
    ram_cell[      36] = 32'h0;  // 32'h6b5d4f25;
    ram_cell[      37] = 32'h0;  // 32'h2ad9cbc0;
    ram_cell[      38] = 32'h0;  // 32'hd5f21b87;
    ram_cell[      39] = 32'h0;  // 32'hb392cc0b;
    ram_cell[      40] = 32'h0;  // 32'haf0300f7;
    ram_cell[      41] = 32'h0;  // 32'h5cc834c5;
    ram_cell[      42] = 32'h0;  // 32'h0e05639f;
    ram_cell[      43] = 32'h0;  // 32'h592e906f;
    ram_cell[      44] = 32'h0;  // 32'h218b1ddb;
    ram_cell[      45] = 32'h0;  // 32'h764485fd;
    ram_cell[      46] = 32'h0;  // 32'hf21d8c7c;
    ram_cell[      47] = 32'h0;  // 32'h9abdd5e1;
    ram_cell[      48] = 32'h0;  // 32'h47e9cccf;
    ram_cell[      49] = 32'h0;  // 32'h2648850f;
    ram_cell[      50] = 32'h0;  // 32'h2277e0ca;
    ram_cell[      51] = 32'h0;  // 32'hfe25401f;
    ram_cell[      52] = 32'h0;  // 32'hbbece3a0;
    ram_cell[      53] = 32'h0;  // 32'h7395561d;
    ram_cell[      54] = 32'h0;  // 32'h57269154;
    ram_cell[      55] = 32'h0;  // 32'h78c77108;
    ram_cell[      56] = 32'h0;  // 32'h53f5f916;
    ram_cell[      57] = 32'h0;  // 32'h130ac35f;
    ram_cell[      58] = 32'h0;  // 32'hb9af1438;
    ram_cell[      59] = 32'h0;  // 32'h16923309;
    ram_cell[      60] = 32'h0;  // 32'h928b159f;
    ram_cell[      61] = 32'h0;  // 32'h2cb3dc2b;
    ram_cell[      62] = 32'h0;  // 32'he3d17939;
    ram_cell[      63] = 32'h0;  // 32'h493845e6;
    ram_cell[      64] = 32'h0;  // 32'h7e146871;
    ram_cell[      65] = 32'h0;  // 32'h2a62579b;
    ram_cell[      66] = 32'h0;  // 32'h54fd857c;
    ram_cell[      67] = 32'h0;  // 32'h899c303c;
    ram_cell[      68] = 32'h0;  // 32'h10e2722f;
    ram_cell[      69] = 32'h0;  // 32'h0553cc2a;
    ram_cell[      70] = 32'h0;  // 32'haecd82bc;
    ram_cell[      71] = 32'h0;  // 32'he6f5e864;
    ram_cell[      72] = 32'h0;  // 32'h164c7841;
    ram_cell[      73] = 32'h0;  // 32'h2db083d5;
    ram_cell[      74] = 32'h0;  // 32'h658e6b7a;
    ram_cell[      75] = 32'h0;  // 32'hec992aac;
    ram_cell[      76] = 32'h0;  // 32'h5d8ab284;
    ram_cell[      77] = 32'h0;  // 32'headdd6b0;
    ram_cell[      78] = 32'h0;  // 32'h392aae3c;
    ram_cell[      79] = 32'h0;  // 32'h6a3c2cb2;
    ram_cell[      80] = 32'h0;  // 32'hc6925b0b;
    ram_cell[      81] = 32'h0;  // 32'h1d417d92;
    ram_cell[      82] = 32'h0;  // 32'hbc198c18;
    ram_cell[      83] = 32'h0;  // 32'h0eb3e021;
    ram_cell[      84] = 32'h0;  // 32'h8f9177db;
    ram_cell[      85] = 32'h0;  // 32'h59455ab5;
    ram_cell[      86] = 32'h0;  // 32'h1e06e6b3;
    ram_cell[      87] = 32'h0;  // 32'h8fbdc3dd;
    ram_cell[      88] = 32'h0;  // 32'h98a263b7;
    ram_cell[      89] = 32'h0;  // 32'h60387cff;
    ram_cell[      90] = 32'h0;  // 32'h43be0c1c;
    ram_cell[      91] = 32'h0;  // 32'h7927cf65;
    ram_cell[      92] = 32'h0;  // 32'h40f15140;
    ram_cell[      93] = 32'h0;  // 32'h97a462c0;
    ram_cell[      94] = 32'h0;  // 32'h19352c8c;
    ram_cell[      95] = 32'h0;  // 32'h5dbfc025;
    ram_cell[      96] = 32'h0;  // 32'he0b3ade2;
    ram_cell[      97] = 32'h0;  // 32'he7b952b7;
    ram_cell[      98] = 32'h0;  // 32'h6fbed911;
    ram_cell[      99] = 32'h0;  // 32'hc534e544;
    ram_cell[     100] = 32'h0;  // 32'h1ac1bb76;
    ram_cell[     101] = 32'h0;  // 32'h14f33970;
    ram_cell[     102] = 32'h0;  // 32'h2d084378;
    ram_cell[     103] = 32'h0;  // 32'h844f021e;
    ram_cell[     104] = 32'h0;  // 32'h7e62caba;
    ram_cell[     105] = 32'h0;  // 32'h9bb69162;
    ram_cell[     106] = 32'h0;  // 32'h44a31c2e;
    ram_cell[     107] = 32'h0;  // 32'hc125417b;
    ram_cell[     108] = 32'h0;  // 32'hfd3dba63;
    ram_cell[     109] = 32'h0;  // 32'h42cf75cb;
    ram_cell[     110] = 32'h0;  // 32'h94be59df;
    ram_cell[     111] = 32'h0;  // 32'h08c31fda;
    ram_cell[     112] = 32'h0;  // 32'h871a9819;
    ram_cell[     113] = 32'h0;  // 32'hb4e2a064;
    ram_cell[     114] = 32'h0;  // 32'h762cea6e;
    ram_cell[     115] = 32'h0;  // 32'hdfc3dcfc;
    ram_cell[     116] = 32'h0;  // 32'h1b499bf9;
    ram_cell[     117] = 32'h0;  // 32'h114afdef;
    ram_cell[     118] = 32'h0;  // 32'hb95c1c2d;
    ram_cell[     119] = 32'h0;  // 32'h22d5385a;
    ram_cell[     120] = 32'h0;  // 32'h37536cd2;
    ram_cell[     121] = 32'h0;  // 32'h4b994e26;
    ram_cell[     122] = 32'h0;  // 32'h4129ab2c;
    ram_cell[     123] = 32'h0;  // 32'hb48df42a;
    ram_cell[     124] = 32'h0;  // 32'h33e9614d;
    ram_cell[     125] = 32'h0;  // 32'h059ce612;
    ram_cell[     126] = 32'h0;  // 32'hffb424d3;
    ram_cell[     127] = 32'h0;  // 32'hdc33d60a;
    ram_cell[     128] = 32'h0;  // 32'h102da57b;
    ram_cell[     129] = 32'h0;  // 32'hec3134e9;
    ram_cell[     130] = 32'h0;  // 32'hb281fb3c;
    ram_cell[     131] = 32'h0;  // 32'h726501c7;
    ram_cell[     132] = 32'h0;  // 32'h785567b6;
    ram_cell[     133] = 32'h0;  // 32'h568fe177;
    ram_cell[     134] = 32'h0;  // 32'hc88656a0;
    ram_cell[     135] = 32'h0;  // 32'ha8e62fb0;
    ram_cell[     136] = 32'h0;  // 32'hc230d402;
    ram_cell[     137] = 32'h0;  // 32'h3b8ff71d;
    ram_cell[     138] = 32'h0;  // 32'h48a39586;
    ram_cell[     139] = 32'h0;  // 32'hc8d2ba46;
    ram_cell[     140] = 32'h0;  // 32'hedab099a;
    ram_cell[     141] = 32'h0;  // 32'h4951d68a;
    ram_cell[     142] = 32'h0;  // 32'h793762d2;
    ram_cell[     143] = 32'h0;  // 32'h2ecad8fa;
    ram_cell[     144] = 32'h0;  // 32'h50ed00d2;
    ram_cell[     145] = 32'h0;  // 32'h07723262;
    ram_cell[     146] = 32'h0;  // 32'h81a73290;
    ram_cell[     147] = 32'h0;  // 32'hed512ed3;
    ram_cell[     148] = 32'h0;  // 32'h85149eea;
    ram_cell[     149] = 32'h0;  // 32'h35bbf9ac;
    ram_cell[     150] = 32'h0;  // 32'h77f8aeca;
    ram_cell[     151] = 32'h0;  // 32'h571cf02b;
    ram_cell[     152] = 32'h0;  // 32'h5b347e2f;
    ram_cell[     153] = 32'h0;  // 32'hd28486ea;
    ram_cell[     154] = 32'h0;  // 32'h8456a44c;
    ram_cell[     155] = 32'h0;  // 32'hd7a3a966;
    ram_cell[     156] = 32'h0;  // 32'h7df32a12;
    ram_cell[     157] = 32'h0;  // 32'h2273943b;
    ram_cell[     158] = 32'h0;  // 32'hc1fedc0f;
    ram_cell[     159] = 32'h0;  // 32'hfe1e40f5;
    ram_cell[     160] = 32'h0;  // 32'ha605c5b4;
    ram_cell[     161] = 32'h0;  // 32'hdad26771;
    ram_cell[     162] = 32'h0;  // 32'h2fdc1b0b;
    ram_cell[     163] = 32'h0;  // 32'h6463dd82;
    ram_cell[     164] = 32'h0;  // 32'h968d72e9;
    ram_cell[     165] = 32'h0;  // 32'h524d0b70;
    ram_cell[     166] = 32'h0;  // 32'h8808f310;
    ram_cell[     167] = 32'h0;  // 32'h0c2655a0;
    ram_cell[     168] = 32'h0;  // 32'h6024b52e;
    ram_cell[     169] = 32'h0;  // 32'h67712a0d;
    ram_cell[     170] = 32'h0;  // 32'h2a52ff36;
    ram_cell[     171] = 32'h0;  // 32'h42579b9b;
    ram_cell[     172] = 32'h0;  // 32'h09617528;
    ram_cell[     173] = 32'h0;  // 32'h550a358d;
    ram_cell[     174] = 32'h0;  // 32'h347b93b9;
    ram_cell[     175] = 32'h0;  // 32'hdc9e145a;
    ram_cell[     176] = 32'h0;  // 32'h30909c3b;
    ram_cell[     177] = 32'h0;  // 32'h308b193c;
    ram_cell[     178] = 32'h0;  // 32'h61f969d6;
    ram_cell[     179] = 32'h0;  // 32'h5b942079;
    ram_cell[     180] = 32'h0;  // 32'haeec9433;
    ram_cell[     181] = 32'h0;  // 32'h9d358ee6;
    ram_cell[     182] = 32'h0;  // 32'hb98f4827;
    ram_cell[     183] = 32'h0;  // 32'h46623a73;
    ram_cell[     184] = 32'h0;  // 32'hb68901a9;
    ram_cell[     185] = 32'h0;  // 32'h735ede6a;
    ram_cell[     186] = 32'h0;  // 32'h00d45e28;
    ram_cell[     187] = 32'h0;  // 32'hc3653ce7;
    ram_cell[     188] = 32'h0;  // 32'hecf45adf;
    ram_cell[     189] = 32'h0;  // 32'h7a7a8e69;
    ram_cell[     190] = 32'h0;  // 32'hf3dfd455;
    ram_cell[     191] = 32'h0;  // 32'h5a780138;
    ram_cell[     192] = 32'h0;  // 32'h96b1ce11;
    ram_cell[     193] = 32'h0;  // 32'h4d1ef516;
    ram_cell[     194] = 32'h0;  // 32'hf7f164fc;
    ram_cell[     195] = 32'h0;  // 32'hd9530c37;
    ram_cell[     196] = 32'h0;  // 32'he298958c;
    ram_cell[     197] = 32'h0;  // 32'hf2edf0c0;
    ram_cell[     198] = 32'h0;  // 32'hd9a5beb8;
    ram_cell[     199] = 32'h0;  // 32'hb00f7369;
    ram_cell[     200] = 32'h0;  // 32'hee4b6442;
    ram_cell[     201] = 32'h0;  // 32'h1c92eb3f;
    ram_cell[     202] = 32'h0;  // 32'hc5a895db;
    ram_cell[     203] = 32'h0;  // 32'h474bad71;
    ram_cell[     204] = 32'h0;  // 32'hd3dfff96;
    ram_cell[     205] = 32'h0;  // 32'h80a550d1;
    ram_cell[     206] = 32'h0;  // 32'h16504033;
    ram_cell[     207] = 32'h0;  // 32'h907d813d;
    ram_cell[     208] = 32'h0;  // 32'hc642410f;
    ram_cell[     209] = 32'h0;  // 32'h735b36bf;
    ram_cell[     210] = 32'h0;  // 32'h7cacce76;
    ram_cell[     211] = 32'h0;  // 32'h6a77eaf7;
    ram_cell[     212] = 32'h0;  // 32'he0508dc4;
    ram_cell[     213] = 32'h0;  // 32'h2c5d241a;
    ram_cell[     214] = 32'h0;  // 32'ha175eea1;
    ram_cell[     215] = 32'h0;  // 32'h5a6fff0a;
    ram_cell[     216] = 32'h0;  // 32'h1b14761a;
    ram_cell[     217] = 32'h0;  // 32'hb325ea8d;
    ram_cell[     218] = 32'h0;  // 32'hb628696c;
    ram_cell[     219] = 32'h0;  // 32'hac6b6895;
    ram_cell[     220] = 32'h0;  // 32'h3628b152;
    ram_cell[     221] = 32'h0;  // 32'h5bf5e20f;
    ram_cell[     222] = 32'h0;  // 32'h39be6774;
    ram_cell[     223] = 32'h0;  // 32'h311def2c;
    ram_cell[     224] = 32'h0;  // 32'hed35b38e;
    ram_cell[     225] = 32'h0;  // 32'h71db03bc;
    ram_cell[     226] = 32'h0;  // 32'h4fcb046c;
    ram_cell[     227] = 32'h0;  // 32'hfd589ea5;
    ram_cell[     228] = 32'h0;  // 32'h43c749a2;
    ram_cell[     229] = 32'h0;  // 32'h6676a8df;
    ram_cell[     230] = 32'h0;  // 32'h0e5556f5;
    ram_cell[     231] = 32'h0;  // 32'ha7dee762;
    ram_cell[     232] = 32'h0;  // 32'h9a16bfcb;
    ram_cell[     233] = 32'h0;  // 32'h523f0307;
    ram_cell[     234] = 32'h0;  // 32'h8655a2f7;
    ram_cell[     235] = 32'h0;  // 32'h2ec156fd;
    ram_cell[     236] = 32'h0;  // 32'hd5618ca1;
    ram_cell[     237] = 32'h0;  // 32'hb69186e6;
    ram_cell[     238] = 32'h0;  // 32'he5ec5352;
    ram_cell[     239] = 32'h0;  // 32'h78a78b72;
    ram_cell[     240] = 32'h0;  // 32'h6a46b9e1;
    ram_cell[     241] = 32'h0;  // 32'h0e385abd;
    ram_cell[     242] = 32'h0;  // 32'h8098722d;
    ram_cell[     243] = 32'h0;  // 32'h9b75b251;
    ram_cell[     244] = 32'h0;  // 32'hd7e74948;
    ram_cell[     245] = 32'h0;  // 32'h11c3bde4;
    ram_cell[     246] = 32'h0;  // 32'h959e76c5;
    ram_cell[     247] = 32'h0;  // 32'h0df6aaba;
    ram_cell[     248] = 32'h0;  // 32'hb3e78a4f;
    ram_cell[     249] = 32'h0;  // 32'hb6d52885;
    ram_cell[     250] = 32'h0;  // 32'h2110a733;
    ram_cell[     251] = 32'h0;  // 32'hc6bd42c5;
    ram_cell[     252] = 32'h0;  // 32'h2434bb3b;
    ram_cell[     253] = 32'h0;  // 32'hfa14a434;
    ram_cell[     254] = 32'h0;  // 32'h9ce80d3f;
    ram_cell[     255] = 32'h0;  // 32'h78053d83;
    // src matrix A
    ram_cell[     256] = 32'h4d2b418a;
    ram_cell[     257] = 32'h34c275b5;
    ram_cell[     258] = 32'h2aefed30;
    ram_cell[     259] = 32'h6d52e82f;
    ram_cell[     260] = 32'h6161d96a;
    ram_cell[     261] = 32'hd07017bb;
    ram_cell[     262] = 32'hfff37878;
    ram_cell[     263] = 32'h53dfb7ce;
    ram_cell[     264] = 32'hd9d0d4aa;
    ram_cell[     265] = 32'h5b9098c5;
    ram_cell[     266] = 32'hd3429622;
    ram_cell[     267] = 32'h656e3436;
    ram_cell[     268] = 32'h9c8f9aae;
    ram_cell[     269] = 32'hbedaf031;
    ram_cell[     270] = 32'ha918bad3;
    ram_cell[     271] = 32'hcb9308a7;
    ram_cell[     272] = 32'h991a7f33;
    ram_cell[     273] = 32'ha65af415;
    ram_cell[     274] = 32'hac5c6847;
    ram_cell[     275] = 32'h48653d8e;
    ram_cell[     276] = 32'h694e328f;
    ram_cell[     277] = 32'h79fa53f6;
    ram_cell[     278] = 32'hff6975d6;
    ram_cell[     279] = 32'hb5ab5ffe;
    ram_cell[     280] = 32'h3d1b1103;
    ram_cell[     281] = 32'hc124eee7;
    ram_cell[     282] = 32'h364ab9de;
    ram_cell[     283] = 32'hebf7b277;
    ram_cell[     284] = 32'h0be03d93;
    ram_cell[     285] = 32'h173b089c;
    ram_cell[     286] = 32'h238a95a3;
    ram_cell[     287] = 32'h790db963;
    ram_cell[     288] = 32'hf89b5228;
    ram_cell[     289] = 32'h7a721901;
    ram_cell[     290] = 32'ha89a4110;
    ram_cell[     291] = 32'hfc8ad06f;
    ram_cell[     292] = 32'h78fcd019;
    ram_cell[     293] = 32'h18eabb22;
    ram_cell[     294] = 32'hc7ad20ba;
    ram_cell[     295] = 32'hbfe2a2f9;
    ram_cell[     296] = 32'h12b0adc6;
    ram_cell[     297] = 32'h0fbf1001;
    ram_cell[     298] = 32'h76f5be60;
    ram_cell[     299] = 32'hfcb69b79;
    ram_cell[     300] = 32'h1f9ae9ef;
    ram_cell[     301] = 32'haf85e749;
    ram_cell[     302] = 32'h58c87f8e;
    ram_cell[     303] = 32'hc1f97479;
    ram_cell[     304] = 32'h99879fb0;
    ram_cell[     305] = 32'hf89bb75e;
    ram_cell[     306] = 32'h5fde99f0;
    ram_cell[     307] = 32'hacb62096;
    ram_cell[     308] = 32'h4c562cde;
    ram_cell[     309] = 32'h671868b6;
    ram_cell[     310] = 32'hc85a3f2c;
    ram_cell[     311] = 32'h6414d3ad;
    ram_cell[     312] = 32'h3ff395b9;
    ram_cell[     313] = 32'h5921f717;
    ram_cell[     314] = 32'h7b5a97b2;
    ram_cell[     315] = 32'hdcf61ede;
    ram_cell[     316] = 32'h56d45c5e;
    ram_cell[     317] = 32'h3bc2075c;
    ram_cell[     318] = 32'h812c8aef;
    ram_cell[     319] = 32'hf1ff51b9;
    ram_cell[     320] = 32'hd19b13eb;
    ram_cell[     321] = 32'h3d7817c4;
    ram_cell[     322] = 32'h30df22c8;
    ram_cell[     323] = 32'h6260a5e5;
    ram_cell[     324] = 32'hc4606963;
    ram_cell[     325] = 32'heb3ed72d;
    ram_cell[     326] = 32'hc65b2221;
    ram_cell[     327] = 32'h24323d82;
    ram_cell[     328] = 32'hff7fe5a8;
    ram_cell[     329] = 32'h07433573;
    ram_cell[     330] = 32'h79e01cad;
    ram_cell[     331] = 32'h86cd5394;
    ram_cell[     332] = 32'hccec8e32;
    ram_cell[     333] = 32'hc5e2d8a2;
    ram_cell[     334] = 32'h2bd5c40c;
    ram_cell[     335] = 32'h8dabdc10;
    ram_cell[     336] = 32'h7de5be4d;
    ram_cell[     337] = 32'hfe676087;
    ram_cell[     338] = 32'h46e8e47c;
    ram_cell[     339] = 32'h4aedf000;
    ram_cell[     340] = 32'hf16f3d35;
    ram_cell[     341] = 32'h342a2ba4;
    ram_cell[     342] = 32'hf6d0f3d7;
    ram_cell[     343] = 32'hbae16bba;
    ram_cell[     344] = 32'h70e891cb;
    ram_cell[     345] = 32'hef755336;
    ram_cell[     346] = 32'hc9cc9dda;
    ram_cell[     347] = 32'h59cede4c;
    ram_cell[     348] = 32'h634411e7;
    ram_cell[     349] = 32'h278eb901;
    ram_cell[     350] = 32'h9f9f5bcd;
    ram_cell[     351] = 32'h8b59be01;
    ram_cell[     352] = 32'hcc88e47d;
    ram_cell[     353] = 32'h4461b28a;
    ram_cell[     354] = 32'hf52cd97e;
    ram_cell[     355] = 32'h20ee0f28;
    ram_cell[     356] = 32'h68f89048;
    ram_cell[     357] = 32'hf26a9752;
    ram_cell[     358] = 32'h613a42d9;
    ram_cell[     359] = 32'h2d5f18d5;
    ram_cell[     360] = 32'h42e094b3;
    ram_cell[     361] = 32'hefc23d00;
    ram_cell[     362] = 32'h0dd294ee;
    ram_cell[     363] = 32'h7bd9391c;
    ram_cell[     364] = 32'h6bb7f285;
    ram_cell[     365] = 32'h390881e5;
    ram_cell[     366] = 32'hc4fccf5b;
    ram_cell[     367] = 32'ha87b4c96;
    ram_cell[     368] = 32'hd2b9acb8;
    ram_cell[     369] = 32'he84e2660;
    ram_cell[     370] = 32'hbee0f170;
    ram_cell[     371] = 32'hffe6bdb2;
    ram_cell[     372] = 32'h095786a1;
    ram_cell[     373] = 32'h06b49fee;
    ram_cell[     374] = 32'h58d31389;
    ram_cell[     375] = 32'h9e2826a5;
    ram_cell[     376] = 32'h60b9c49d;
    ram_cell[     377] = 32'hef1eaeae;
    ram_cell[     378] = 32'h59a7b87b;
    ram_cell[     379] = 32'hd5260cfa;
    ram_cell[     380] = 32'hc8449d42;
    ram_cell[     381] = 32'h796b246b;
    ram_cell[     382] = 32'h0a13bd90;
    ram_cell[     383] = 32'h0a7e2a7e;
    ram_cell[     384] = 32'h8acaf855;
    ram_cell[     385] = 32'h0d466814;
    ram_cell[     386] = 32'h0b0a162e;
    ram_cell[     387] = 32'h95593387;
    ram_cell[     388] = 32'h6f2460af;
    ram_cell[     389] = 32'hfc040da9;
    ram_cell[     390] = 32'h52f38164;
    ram_cell[     391] = 32'h406ee0cc;
    ram_cell[     392] = 32'h47b969aa;
    ram_cell[     393] = 32'h196574e0;
    ram_cell[     394] = 32'h9fd61645;
    ram_cell[     395] = 32'hb10b0f3d;
    ram_cell[     396] = 32'he600106b;
    ram_cell[     397] = 32'hf560cadf;
    ram_cell[     398] = 32'h2148b11b;
    ram_cell[     399] = 32'h6c178f12;
    ram_cell[     400] = 32'he4f1b976;
    ram_cell[     401] = 32'hb2b7bc75;
    ram_cell[     402] = 32'he98a3b2b;
    ram_cell[     403] = 32'h7713b46d;
    ram_cell[     404] = 32'hd1ed2909;
    ram_cell[     405] = 32'h7679c5fc;
    ram_cell[     406] = 32'h120d3536;
    ram_cell[     407] = 32'h5fdfaaca;
    ram_cell[     408] = 32'hd244cef6;
    ram_cell[     409] = 32'ha0ead1d4;
    ram_cell[     410] = 32'h1d1feebf;
    ram_cell[     411] = 32'he6720564;
    ram_cell[     412] = 32'he0d03557;
    ram_cell[     413] = 32'h914d17cc;
    ram_cell[     414] = 32'hcefbeb2b;
    ram_cell[     415] = 32'h2800c446;
    ram_cell[     416] = 32'h2e4b7310;
    ram_cell[     417] = 32'hbd680ca0;
    ram_cell[     418] = 32'h934e21f4;
    ram_cell[     419] = 32'he093ce7a;
    ram_cell[     420] = 32'h9310464d;
    ram_cell[     421] = 32'h4db0d1b2;
    ram_cell[     422] = 32'h278288a8;
    ram_cell[     423] = 32'hcf92c8ec;
    ram_cell[     424] = 32'hef725351;
    ram_cell[     425] = 32'hf072e7f3;
    ram_cell[     426] = 32'h8babcc8c;
    ram_cell[     427] = 32'h83233b4e;
    ram_cell[     428] = 32'hfb40c3ad;
    ram_cell[     429] = 32'hc5fca635;
    ram_cell[     430] = 32'ha0be4240;
    ram_cell[     431] = 32'h61331265;
    ram_cell[     432] = 32'h9acfc335;
    ram_cell[     433] = 32'hf61ec2e0;
    ram_cell[     434] = 32'h184d89e0;
    ram_cell[     435] = 32'heb4bc9fe;
    ram_cell[     436] = 32'h26d67441;
    ram_cell[     437] = 32'haaa8090a;
    ram_cell[     438] = 32'h3f7a730e;
    ram_cell[     439] = 32'he9effde2;
    ram_cell[     440] = 32'h75bd1ce4;
    ram_cell[     441] = 32'h2887fb98;
    ram_cell[     442] = 32'h263f7d77;
    ram_cell[     443] = 32'h639ebb84;
    ram_cell[     444] = 32'hbd902179;
    ram_cell[     445] = 32'hb3e6f2e1;
    ram_cell[     446] = 32'h988f0077;
    ram_cell[     447] = 32'h31ae11f1;
    ram_cell[     448] = 32'h443e9caa;
    ram_cell[     449] = 32'h7faaac30;
    ram_cell[     450] = 32'h6243ac86;
    ram_cell[     451] = 32'h094b44a5;
    ram_cell[     452] = 32'h4d552e51;
    ram_cell[     453] = 32'h59e2d9ca;
    ram_cell[     454] = 32'hb84d5116;
    ram_cell[     455] = 32'h1de2ec7e;
    ram_cell[     456] = 32'h98a8d767;
    ram_cell[     457] = 32'he7b75327;
    ram_cell[     458] = 32'he9579f8d;
    ram_cell[     459] = 32'h767eeded;
    ram_cell[     460] = 32'h837412c8;
    ram_cell[     461] = 32'ha9743fd7;
    ram_cell[     462] = 32'h12d853c1;
    ram_cell[     463] = 32'h4ff86093;
    ram_cell[     464] = 32'h776a6cb0;
    ram_cell[     465] = 32'h32f6f0dc;
    ram_cell[     466] = 32'h39c09aca;
    ram_cell[     467] = 32'hda030962;
    ram_cell[     468] = 32'h73dec5b5;
    ram_cell[     469] = 32'hba279e94;
    ram_cell[     470] = 32'had249a48;
    ram_cell[     471] = 32'hae3ad2b7;
    ram_cell[     472] = 32'h2f90fad8;
    ram_cell[     473] = 32'hf343d4dc;
    ram_cell[     474] = 32'h3d6069be;
    ram_cell[     475] = 32'h4f27787c;
    ram_cell[     476] = 32'h4750dbb3;
    ram_cell[     477] = 32'h4a22622d;
    ram_cell[     478] = 32'h8ebf86a5;
    ram_cell[     479] = 32'hda119b95;
    ram_cell[     480] = 32'h82248791;
    ram_cell[     481] = 32'ha9514715;
    ram_cell[     482] = 32'ha5280f84;
    ram_cell[     483] = 32'h024044cd;
    ram_cell[     484] = 32'hcee9b099;
    ram_cell[     485] = 32'h71fdb416;
    ram_cell[     486] = 32'h3fd7b24d;
    ram_cell[     487] = 32'hdc69452a;
    ram_cell[     488] = 32'hd3aa15ea;
    ram_cell[     489] = 32'h125ad86f;
    ram_cell[     490] = 32'ha06ff6c0;
    ram_cell[     491] = 32'hd6c39fdf;
    ram_cell[     492] = 32'h5397b6d2;
    ram_cell[     493] = 32'h137ba6b5;
    ram_cell[     494] = 32'h1a32284e;
    ram_cell[     495] = 32'h57731f21;
    ram_cell[     496] = 32'hdd5fe890;
    ram_cell[     497] = 32'he2df7d7a;
    ram_cell[     498] = 32'h129b7efc;
    ram_cell[     499] = 32'h3731ed5e;
    ram_cell[     500] = 32'h05108a7a;
    ram_cell[     501] = 32'h8872f3e5;
    ram_cell[     502] = 32'hd05418e6;
    ram_cell[     503] = 32'h8c8ed2ad;
    ram_cell[     504] = 32'hf71dc447;
    ram_cell[     505] = 32'h3fab09ab;
    ram_cell[     506] = 32'h323201c0;
    ram_cell[     507] = 32'he9c20715;
    ram_cell[     508] = 32'h1800ca85;
    ram_cell[     509] = 32'ha0d293e5;
    ram_cell[     510] = 32'h6bb8581a;
    ram_cell[     511] = 32'h337a9086;
    // src matrix B
    ram_cell[     512] = 32'hc8ffbf74;
    ram_cell[     513] = 32'he7cb2a86;
    ram_cell[     514] = 32'h47e4620a;
    ram_cell[     515] = 32'h5d075b09;
    ram_cell[     516] = 32'hfe61f95e;
    ram_cell[     517] = 32'h01739c0f;
    ram_cell[     518] = 32'h1334b90d;
    ram_cell[     519] = 32'hc69285da;
    ram_cell[     520] = 32'hd76dd3b9;
    ram_cell[     521] = 32'hf1f99cc5;
    ram_cell[     522] = 32'ha92ff748;
    ram_cell[     523] = 32'hd7ad269c;
    ram_cell[     524] = 32'h9805ebb4;
    ram_cell[     525] = 32'h26a17a35;
    ram_cell[     526] = 32'h8d716e65;
    ram_cell[     527] = 32'h12b5bca9;
    ram_cell[     528] = 32'h11f0d599;
    ram_cell[     529] = 32'he5e2e9e5;
    ram_cell[     530] = 32'h0bf60f3d;
    ram_cell[     531] = 32'hdc47148e;
    ram_cell[     532] = 32'h94af1319;
    ram_cell[     533] = 32'h843befa2;
    ram_cell[     534] = 32'h4dc473fd;
    ram_cell[     535] = 32'h25c51761;
    ram_cell[     536] = 32'h13f96eef;
    ram_cell[     537] = 32'h382d63e1;
    ram_cell[     538] = 32'hb8a9dbd8;
    ram_cell[     539] = 32'h1f377ef0;
    ram_cell[     540] = 32'h9c48fa10;
    ram_cell[     541] = 32'hbb850d46;
    ram_cell[     542] = 32'h5a9fcd17;
    ram_cell[     543] = 32'h8ccc9f30;
    ram_cell[     544] = 32'he63420e7;
    ram_cell[     545] = 32'h423a098c;
    ram_cell[     546] = 32'hdd9fcdfb;
    ram_cell[     547] = 32'hfe451d7e;
    ram_cell[     548] = 32'h9f59a2a9;
    ram_cell[     549] = 32'h9ab84fa9;
    ram_cell[     550] = 32'hbd30ad2a;
    ram_cell[     551] = 32'h65f763d1;
    ram_cell[     552] = 32'heb026587;
    ram_cell[     553] = 32'h2ff1e366;
    ram_cell[     554] = 32'hae78e8c1;
    ram_cell[     555] = 32'h807f3981;
    ram_cell[     556] = 32'h8de1576a;
    ram_cell[     557] = 32'h4a7ee197;
    ram_cell[     558] = 32'h6c9d5c0e;
    ram_cell[     559] = 32'h2c5a0ed2;
    ram_cell[     560] = 32'h003bc89d;
    ram_cell[     561] = 32'haa2b99fc;
    ram_cell[     562] = 32'hf001be07;
    ram_cell[     563] = 32'h4574d264;
    ram_cell[     564] = 32'heee811d5;
    ram_cell[     565] = 32'hf770edcd;
    ram_cell[     566] = 32'h4df5b74f;
    ram_cell[     567] = 32'he0addbed;
    ram_cell[     568] = 32'hec296050;
    ram_cell[     569] = 32'hefbf1450;
    ram_cell[     570] = 32'h01ddaf3f;
    ram_cell[     571] = 32'haf1b0cfe;
    ram_cell[     572] = 32'h829e2de2;
    ram_cell[     573] = 32'hceaf9ec4;
    ram_cell[     574] = 32'h7c39462f;
    ram_cell[     575] = 32'hca5a19ca;
    ram_cell[     576] = 32'h1825dfaf;
    ram_cell[     577] = 32'h14b93aab;
    ram_cell[     578] = 32'hdd5f65a9;
    ram_cell[     579] = 32'h32225aba;
    ram_cell[     580] = 32'hd501c8df;
    ram_cell[     581] = 32'h7507d2b2;
    ram_cell[     582] = 32'hc8391c09;
    ram_cell[     583] = 32'h81455d0b;
    ram_cell[     584] = 32'hbb05a145;
    ram_cell[     585] = 32'haffa2e0a;
    ram_cell[     586] = 32'hc09871f0;
    ram_cell[     587] = 32'h6137caa0;
    ram_cell[     588] = 32'h8d48776b;
    ram_cell[     589] = 32'hfa9cb061;
    ram_cell[     590] = 32'h4cfe396e;
    ram_cell[     591] = 32'h3a18dddc;
    ram_cell[     592] = 32'h213471a3;
    ram_cell[     593] = 32'hc8af036f;
    ram_cell[     594] = 32'hd32b9f48;
    ram_cell[     595] = 32'h9a25bca4;
    ram_cell[     596] = 32'h1558fed9;
    ram_cell[     597] = 32'h917a116c;
    ram_cell[     598] = 32'h9f8a11c5;
    ram_cell[     599] = 32'h536b3b93;
    ram_cell[     600] = 32'h327d7b91;
    ram_cell[     601] = 32'h007e337b;
    ram_cell[     602] = 32'h1c05f269;
    ram_cell[     603] = 32'he15a2bb5;
    ram_cell[     604] = 32'h17ca14f7;
    ram_cell[     605] = 32'h640bcf67;
    ram_cell[     606] = 32'h9b101ada;
    ram_cell[     607] = 32'h49bf3176;
    ram_cell[     608] = 32'h3bfd9b1e;
    ram_cell[     609] = 32'hff58539c;
    ram_cell[     610] = 32'hcb28ffb2;
    ram_cell[     611] = 32'h3635ed75;
    ram_cell[     612] = 32'h70610386;
    ram_cell[     613] = 32'h1a04284e;
    ram_cell[     614] = 32'h3bbb4f77;
    ram_cell[     615] = 32'h00a32658;
    ram_cell[     616] = 32'hc073661d;
    ram_cell[     617] = 32'hd03ffa14;
    ram_cell[     618] = 32'h63e5154a;
    ram_cell[     619] = 32'ha11ba8e3;
    ram_cell[     620] = 32'h1863cf54;
    ram_cell[     621] = 32'h69d53d99;
    ram_cell[     622] = 32'h4358ea1d;
    ram_cell[     623] = 32'h1fe33379;
    ram_cell[     624] = 32'h40c068c3;
    ram_cell[     625] = 32'h40c6a89e;
    ram_cell[     626] = 32'h3d18abb6;
    ram_cell[     627] = 32'h67d2cdaf;
    ram_cell[     628] = 32'ha23c4d70;
    ram_cell[     629] = 32'h64bb6fee;
    ram_cell[     630] = 32'hcec78b3e;
    ram_cell[     631] = 32'h10f84227;
    ram_cell[     632] = 32'h42fb7e77;
    ram_cell[     633] = 32'h9a9d1dbb;
    ram_cell[     634] = 32'h9e4044ac;
    ram_cell[     635] = 32'h0b8f86a1;
    ram_cell[     636] = 32'hc1132f6b;
    ram_cell[     637] = 32'h055feefd;
    ram_cell[     638] = 32'hc3b75284;
    ram_cell[     639] = 32'hb53be575;
    ram_cell[     640] = 32'h17380e04;
    ram_cell[     641] = 32'hea182d36;
    ram_cell[     642] = 32'h0dbee6b9;
    ram_cell[     643] = 32'hb177bee5;
    ram_cell[     644] = 32'h425058a0;
    ram_cell[     645] = 32'h8679a596;
    ram_cell[     646] = 32'hb1542763;
    ram_cell[     647] = 32'h89a483ab;
    ram_cell[     648] = 32'h3713441b;
    ram_cell[     649] = 32'h5b92a31f;
    ram_cell[     650] = 32'h44495938;
    ram_cell[     651] = 32'ha21c0f02;
    ram_cell[     652] = 32'hc5bbfad5;
    ram_cell[     653] = 32'h74d506cc;
    ram_cell[     654] = 32'h1e9a3271;
    ram_cell[     655] = 32'h292e1c64;
    ram_cell[     656] = 32'hc0f6ea31;
    ram_cell[     657] = 32'h4f6b9c20;
    ram_cell[     658] = 32'hfbe03e7a;
    ram_cell[     659] = 32'h5c198900;
    ram_cell[     660] = 32'h253c9845;
    ram_cell[     661] = 32'h414845d9;
    ram_cell[     662] = 32'h41a588ba;
    ram_cell[     663] = 32'h35766109;
    ram_cell[     664] = 32'h6dc2af94;
    ram_cell[     665] = 32'h138c4144;
    ram_cell[     666] = 32'h5e9dea50;
    ram_cell[     667] = 32'hc99e83b3;
    ram_cell[     668] = 32'he248a3d6;
    ram_cell[     669] = 32'hea12cb34;
    ram_cell[     670] = 32'h2369c6b3;
    ram_cell[     671] = 32'h3e915684;
    ram_cell[     672] = 32'h0a97a353;
    ram_cell[     673] = 32'h51a9e7f9;
    ram_cell[     674] = 32'h97c80d44;
    ram_cell[     675] = 32'ha0769e28;
    ram_cell[     676] = 32'h0f6a0db9;
    ram_cell[     677] = 32'h24d6e955;
    ram_cell[     678] = 32'he912835f;
    ram_cell[     679] = 32'h99bad5ea;
    ram_cell[     680] = 32'h1e6b7fcd;
    ram_cell[     681] = 32'ha2148881;
    ram_cell[     682] = 32'hb792db74;
    ram_cell[     683] = 32'h746463ab;
    ram_cell[     684] = 32'hb29e0f24;
    ram_cell[     685] = 32'h129d9302;
    ram_cell[     686] = 32'h2930505c;
    ram_cell[     687] = 32'h8e2a7d22;
    ram_cell[     688] = 32'hbe4716d0;
    ram_cell[     689] = 32'h42c74ef5;
    ram_cell[     690] = 32'h935c9e0c;
    ram_cell[     691] = 32'hbeed486c;
    ram_cell[     692] = 32'h7597224c;
    ram_cell[     693] = 32'hf6fabc1b;
    ram_cell[     694] = 32'hf8242d4c;
    ram_cell[     695] = 32'h7b37348b;
    ram_cell[     696] = 32'hda8d4082;
    ram_cell[     697] = 32'h83e80d59;
    ram_cell[     698] = 32'haffda08c;
    ram_cell[     699] = 32'h65665335;
    ram_cell[     700] = 32'h00fa9dcf;
    ram_cell[     701] = 32'he1094c4d;
    ram_cell[     702] = 32'haf1b7d80;
    ram_cell[     703] = 32'ha323749e;
    ram_cell[     704] = 32'h5ddc0f92;
    ram_cell[     705] = 32'h9cf8eadb;
    ram_cell[     706] = 32'h62f419f6;
    ram_cell[     707] = 32'h8c658d30;
    ram_cell[     708] = 32'h78f811e5;
    ram_cell[     709] = 32'hb274c7ce;
    ram_cell[     710] = 32'hdeadbe92;
    ram_cell[     711] = 32'h7667552e;
    ram_cell[     712] = 32'hd9ff3567;
    ram_cell[     713] = 32'h5fc66b5a;
    ram_cell[     714] = 32'h6813b5f6;
    ram_cell[     715] = 32'hcfcf6f2e;
    ram_cell[     716] = 32'h1631c125;
    ram_cell[     717] = 32'hed15bc9e;
    ram_cell[     718] = 32'h25374fe2;
    ram_cell[     719] = 32'h79c5ce48;
    ram_cell[     720] = 32'hd5bc90e2;
    ram_cell[     721] = 32'h35cd59d0;
    ram_cell[     722] = 32'he4fdacd6;
    ram_cell[     723] = 32'h1c7bb44f;
    ram_cell[     724] = 32'h4864dbd3;
    ram_cell[     725] = 32'hc5b728d6;
    ram_cell[     726] = 32'h5bd0c145;
    ram_cell[     727] = 32'hc96f33f1;
    ram_cell[     728] = 32'h3b9f62dd;
    ram_cell[     729] = 32'ha9406139;
    ram_cell[     730] = 32'h97bde67e;
    ram_cell[     731] = 32'h48bbc35d;
    ram_cell[     732] = 32'h28d27cd4;
    ram_cell[     733] = 32'h34ffe427;
    ram_cell[     734] = 32'h049c31b3;
    ram_cell[     735] = 32'hed2c6d20;
    ram_cell[     736] = 32'h21fb5071;
    ram_cell[     737] = 32'hfd8bbc98;
    ram_cell[     738] = 32'h84930252;
    ram_cell[     739] = 32'h98d6660d;
    ram_cell[     740] = 32'hedf716dc;
    ram_cell[     741] = 32'h76fad51b;
    ram_cell[     742] = 32'h275c4b66;
    ram_cell[     743] = 32'hc7bb01cf;
    ram_cell[     744] = 32'h7e1c222a;
    ram_cell[     745] = 32'hdcd611de;
    ram_cell[     746] = 32'ha840c990;
    ram_cell[     747] = 32'h58da43fa;
    ram_cell[     748] = 32'hb890965a;
    ram_cell[     749] = 32'haa870b41;
    ram_cell[     750] = 32'hbc1df05f;
    ram_cell[     751] = 32'hfbf524a1;
    ram_cell[     752] = 32'h9df9c7f2;
    ram_cell[     753] = 32'hcef9950b;
    ram_cell[     754] = 32'hb149eda9;
    ram_cell[     755] = 32'h634a1d1a;
    ram_cell[     756] = 32'hec76e3b1;
    ram_cell[     757] = 32'h39ca7a55;
    ram_cell[     758] = 32'h13aee2a9;
    ram_cell[     759] = 32'h4b2bf25a;
    ram_cell[     760] = 32'h95724088;
    ram_cell[     761] = 32'hf6d5fb57;
    ram_cell[     762] = 32'hf506c872;
    ram_cell[     763] = 32'h3c383443;
    ram_cell[     764] = 32'h40f9769f;
    ram_cell[     765] = 32'h6a67453f;
    ram_cell[     766] = 32'h6c1fd01a;
    ram_cell[     767] = 32'he60b21b8;
end

endmodule

